module shift_counter (in, login, out);
   //We assume that maximum value of n is 32, so log(32) is 5, so we maximum use 5-bit register. so range is 0-5 bit.
   input in;
   input logg;

   input [6:0] in;
   input [6:0] login;
   output out;
   
   output 
   
   
endmodule